// 32-bit representation

W4_0 = 32'b 0111 1111 1111 1111 0000 0000 0000 0000;

W4_1 = 32'b 0000 0000 0000 0000 1000 0000 0000 0000;

W4_2 = 32'b 1000 0000 0000 0000 0000 0000 0000 0000; // W4_2 = -W4_0

W4_3 = 32'b 0000 0000 0000 0000 0111 1111 1111 1111; // W4_3 = -W4_1



// 1 / sqrt(2) times 2e15 in binary 16bit is 0101 1010 1000 0010

// -1 / sqrt(2) times 2e15 in binary 16bit is 1010 0101 0111 1110


W8_0 = 32'b 0111 1111 1111 1111 0000 0000 0000 0000;

W8_1 = 32'b 0101 1010 1000 0010 1010 0101 0111 1110;

W8_2 = 32'b 0000 0000 0000 0000 1000 0000 0000 0000;

W8_3 = 32'b 1010 0101 0111 1110 1010 0101 0111 1110;

W8_4 = 32'b 1000 0000 0000 0000 0000 0000 0000 0000; // W8_4 = -W8_0

W8_5 = 32'b 1010 0101 0111 1110 0101 1010 1000 0010; // W8_5 = -W8_1

W8_6 = 32'b 0000 0000 0000 0000 0111 1111 1111 1111; // W8_6 = -W8_2

W8_7 = 32'b 0101 1010 1000 0010 0101 1010 1000 0010; // W8_7 = -W8_3